magic
tech sky130A
timestamp 1712357396
<< nwell >>
rect -400 -100 -100 300
<< nmos >>
rect -260 -300 -245 -200
<< pmos >>
rect -260 -55 -245 155
<< ndiff >>
rect -300 -210 -260 -200
rect -300 -290 -295 -210
rect -270 -290 -260 -210
rect -300 -300 -260 -290
rect -245 -210 -200 -200
rect -245 -290 -235 -210
rect -205 -290 -200 -210
rect -245 -300 -200 -290
<< pdiff >>
rect -315 145 -260 155
rect -315 -45 -305 145
rect -270 -45 -260 145
rect -315 -55 -260 -45
rect -245 145 -190 155
rect -245 -45 -235 145
rect -195 -45 -190 145
rect -245 -55 -190 -45
<< ndiffc >>
rect -295 -290 -270 -210
rect -235 -290 -205 -210
<< pdiffc >>
rect -305 -45 -270 145
rect -235 -45 -195 145
<< psubdiff >>
rect -305 -345 -195 -330
rect -305 -375 -290 -345
rect -210 -375 -195 -345
rect -305 -390 -195 -375
<< nsubdiff >>
rect -330 260 -165 275
rect -330 230 -315 260
rect -180 230 -165 260
rect -330 215 -165 230
<< psubdiffcont >>
rect -290 -375 -210 -345
<< nsubdiffcont >>
rect -315 230 -180 260
<< poly >>
rect -260 155 -245 175
rect -260 -125 -245 -55
rect -325 -130 -245 -125
rect -325 -155 -310 -130
rect -285 -155 -245 -130
rect -325 -160 -245 -155
rect -210 -130 -170 -125
rect -210 -150 -200 -130
rect -180 -150 -170 -130
rect -210 -160 -170 -150
rect -260 -200 -245 -160
rect -260 -315 -245 -300
<< polycont >>
rect -310 -155 -285 -130
rect -200 -150 -180 -130
<< locali >>
rect -330 270 -165 275
rect -330 260 -300 270
rect -210 260 -165 270
rect -330 230 -315 260
rect -180 230 -165 260
rect -330 220 -300 230
rect -210 220 -165 230
rect -330 215 -165 220
rect -310 155 -270 215
rect -315 145 -265 155
rect -315 -45 -305 145
rect -270 -45 -265 145
rect -315 -55 -265 -45
rect -240 145 -190 155
rect -240 -45 -235 145
rect -195 -45 -190 145
rect -240 -55 -190 -45
rect -240 -125 -200 -55
rect -325 -130 -275 -125
rect -325 -155 -310 -130
rect -285 -155 -275 -130
rect -325 -160 -275 -155
rect -240 -130 -170 -125
rect -240 -150 -200 -130
rect -180 -150 -170 -130
rect -240 -160 -170 -150
rect -300 -210 -265 -200
rect -300 -290 -295 -210
rect -270 -290 -265 -210
rect -300 -300 -265 -290
rect -240 -210 -200 -160
rect -240 -290 -235 -210
rect -205 -290 -200 -210
rect -240 -300 -200 -290
rect -300 -335 -270 -300
rect -300 -340 -200 -335
rect -300 -345 -280 -340
rect -220 -345 -200 -340
rect -300 -375 -290 -345
rect -210 -375 -200 -345
rect -300 -380 -280 -375
rect -220 -380 -200 -375
rect -300 -385 -200 -380
<< viali >>
rect -300 260 -210 270
rect -300 230 -210 260
rect -300 220 -210 230
rect -310 -155 -285 -130
rect -200 -150 -180 -130
rect -280 -345 -220 -340
rect -280 -375 -220 -345
rect -280 -380 -220 -375
<< metal1 >>
rect -730 270 285 275
rect -730 220 -300 270
rect -210 220 285 270
rect -730 215 285 220
rect -415 -130 -275 -125
rect -415 -155 -310 -130
rect -285 -155 -275 -130
rect -415 -160 -275 -155
rect -240 -130 10 -125
rect -240 -150 -200 -130
rect -180 -150 10 -130
rect -240 -160 10 -150
rect -735 -340 280 -330
rect -735 -380 -280 -340
rect -220 -380 280 -340
rect -735 -390 280 -380
<< labels >>
rlabel metal1 170 240 170 240 1 vdd
rlabel metal1 190 -360 190 -360 1 vss
rlabel metal1 -10 -150 5 -135 1 out
rlabel metal1 -410 -150 -395 -135 1 in
<< end >>
